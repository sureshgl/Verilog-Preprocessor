/* jjjhbjmnb
jhbhjbhjkbmnbhjb 
bhjbknmnbjkb */
module undef_testData;
using beforing undoing third_defination
using beforing undoing second_defination

endmodule
