module ifdef_elseif_else_end_testData();

initial
begin

	$display(" TYPE_1 message ");
	abc_type_1
end

begin
$display(" TYPE_8 message ");
	module ifdef_in_statement_else();
endmodule;
end

type2
    tmp_data[8:0] = {write_data[8:0]}
    tmp = abcccc;

entered else in type_3


assign power = (VDD_buf=== 1'b1 && VSS_buf=== 1'b0) ? 1:0;

always @(VDD_buf or VSS_buf )
begin // {
        if(VDD_buf !== 1'b1) begin // {
                uut.task_corrupt_memory_x;
                uut.task_corrupt_output_x;
                if( MES_CNTRL >= ERROR )
                begin // {
                  $display("<<LSI_MEM_111HS_ERROR: VDD is invalid. Corrupting Memory & output>> at time=%t; instance=%m\n",$realtime);
                end // }
        end // }
        if(VSS_buf !== 1'b0) begin // {
                uut.task_corrupt_memory_x;
                uut.task_corrupt_output_x;
                if( MES_CNTRL >= ERROR )
                begin // {
                  $display("<<LSI_MEM_111HS_ERROR: VSS is invalid. Corrupting Memory & output>> at time=%t; instance=%m\n",$realtime);
                end // }
        end // }
end     // }




in ifndef type6


begin
	in else of ifndef TYPE_5


tmp_data= 1111;
                 tmp_data = 7777777;

begin
    tmp_data[43:0] =ABC;
                tmp_data = 555;

endmodule