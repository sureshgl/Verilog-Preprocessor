/* jjjhbjmnb
jhbhjbhjkbmnbhjb 
bhjbknmnbjkb */
module undef_testData;
`define one first_defination
`define two second_defination
`define three third_defination
using beforing undoing `three
using beforing undoing `two
`undef three
`undef two
// undoingggggggg
endmodule