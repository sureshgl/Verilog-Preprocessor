module reset_all_testData;
using the defination before reset second_defination
using the defination before reset
endmodule;