//define rule shud end with newline
module xyz;
******************
shouldnot process this xyz
endmodule

module define_rule_testdata;
abc abc ;
xyz xyz ;

result = 5 + 5;   5   $display("Inside ADD5 macro. Scope is %m");
2 + 2
"Hello world!"
20
1
1vg@#|1
1
2+1+2+2
32'h0076f020
5
endmodule

module abc;
******************
shouldnot process this
endmodule