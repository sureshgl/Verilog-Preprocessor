module reset_all_testData;
`define one first_defination
`define two second_defination
`define three third_defination
using the defination before reset `two
`resetall
using the defination before reset
endmodule;