module search_path_testData;
`define search searching_in_search_path
in search_path_test;

`search
endmodule