 some text before instantiation_testData;
 abc abc ;
 xyz xyz ;
 
 module instantiation_testData;
 some text inside instantiation_testData;
 
 
 
 instantiation_part2_GWQAUSSR#(.a(12),.b(34)) nameofinstance (); 
 
 processing next **********;
 
 
 second_declaration_XDYFQXHV#() second(); 
 
 
 
endmodule


some text before instantiation_testData;
abc abc ;
xyz xyz ;

module instantiation_testData;
	some text inside instantiation_testData;

	
	instantiation_part2_GVUBMZOF#(.a(12),.b(34)) nameofinstance ();

	processing next **********;
	
	second_declaration_PVTCLXVX#() second();

	`in_second;

endmodule

